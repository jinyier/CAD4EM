`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:38:16 02/05/2020
// Design Name:   aes_192
// Module Name:   D:/TestData/aspdac_tool/aes_cep/aes_cep/aes_top/aes_192/tb.v
// Project Name:  aes_192
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: aes_192
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	reg clk;
	reg rst;
	reg start;
	reg [127:0] state;
	reg [191:0] key;
	// Outputs
	wire out1;
	wire kf1;
	wire out_valid;

	// Instantiate the Unit Under Test (UUT)
	aes_192 uut (
		.clk(clk), 
		.rst(rst), 
		.start(start), 
		.state(state), 
		.key(key),
		.out1(out1), 
		.kf1(kf1),
		.out_valid(out_valid)
	);

  parameter CLK_HALF_PERIOD = 10;
  parameter CLK_PERIOD = 2 * CLK_HALF_PERIOD;
  parameter CLK_SAMPLE_HALF_PERIOD = 5;
   reg			sample_clk;
 
   always
    begin : clk_gen
      #CLK_HALF_PERIOD;
      clk = !clk;
    end // clk_gen

	
	  always
    begin : sample_clk_gen
      #CLK_SAMPLE_HALF_PERIOD;
      sample_clk = !sample_clk;
    end // sample_clk_gen

  task init_sim;
    begin

      clk     = 0;
      rst = 1;
      sample_clk=0;
      start=0;
      key = 128'hffffffffffffffffffffffffffffffff;
      state  = 128'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa;
    end
  endtask // init_sim

  task reset_dut;
    begin
      rst = 1;
      #(2 * CLK_PERIOD);
      rst = 0;
    end
  endtask // reset_dut

initial $readmemh("semi_plain.txt", ktp_data);


	integer i=0;
	parameter num=1000;
	reg [255:0] ktp_data [num:1];

initial	
   begin : main
      $display("   -= Testbench for AES started =-");
      $display("    ==============================");
      $display("");

      init_sim();
		reset_dut();
 
	for(i=1;i<=num;i=i+1)
	begin
	  key = ktp_data[i][255:128];
      state = ktp_data[i][127:0];
      start=1;
      #(2 * CLK_PERIOD); 
      start=0;
	  #(26 * CLK_PERIOD); 	
	end
      //display_test_results();
        //#(100 * CLK_PERIOD);
      $display("");
      $display("*** AES simulation done. ***");
      $finish;
    end // main
	 
    reg [1407:0] data1,data2;
		always@(posedge clk)
		
		begin
			if(rst)
    data1<= 0;
			else
			data1<={uut.s1[43],uut.s6[105],uut.s4[107],uut.s3[10],uut.s11[70],uut.s2[88],uut.s2[43],uut.s7[68],uut.s9[110],uut.s1[52],uut.s3[9],uut.s1[62],uut.s2[62],uut.s6[46],uut.s6[18],uut.s8[6],uut.s2[33],uut.s2[52],uut.s5[117],uut.s9[88],uut.s9[34],uut.s11[90],uut.s8[124],uut.s4[113],uut.s2[70],uut.s10[44],uut.s5[19],uut.s1[108],uut.s8[91],uut.s7[101],uut.s9[13],uut.s9[67],uut.s6[1],uut.s5[43],uut.s7[60],uut.s4[43],uut.s11[106],uut.s1[15],uut.s4[112],uut.s6[75],uut.s1[111],uut.s3[82],uut.s7[78],uut.s4[69],uut.s3[25],uut.s6[122],uut.s9[40],uut.s5[68],uut.s9[55],uut.s7[52],uut.s5[87],uut.s5[92],uut.s8[0],uut.s9[62],uut.s5[122],uut.s11[77],uut.s11[75],uut.s1[33],uut.s1[38],uut.s4[125],uut.s9[69],uut.s4[53],uut.s10[96],uut.s6[94],uut.s1[56],uut.s3[16],uut.s10[21],uut.s5[61],uut.s8[21],uut.s2[126],uut.s2[27],uut.s1[82],uut.s8[71],uut.s9[49],uut.s4[111],uut.s3[18],uut.s8[1],uut.s9[115],uut.s7[67],uut.s8[54],uut.s9[98],uut.s11[107],uut.s6[55],uut.s1[90],uut.s11[44],uut.s8[32],uut.s9[87],uut.s8[83],uut.s11[108],uut.s5[25],uut.s10[40],uut.s1[54],uut.s8[67],uut.s7[25],uut.s4[118],uut.s9[104],uut.s3[96],uut.s8[96],uut.s3[86],uut.s2[96],uut.s11[104],uut.s10[100],uut.s6[78],uut.s2[31],uut.s3[75],uut.s2[90],uut.s5[34],uut.s9[116],uut.s1[41],uut.s3[59],uut.s10[28],uut.s9[57],uut.s6[109],uut.s4[61],uut.s11[33],uut.s6[101],uut.s8[78],uut.s10[38],uut.s9[76],uut.s9[81],uut.s11[126],uut.s1[39],uut.s8[88],uut.s7[89],uut.s7[47],uut.s8[109],uut.s8[19],uut.s11[32],uut.s2[24],uut.s4[101],uut.s7[66],uut.s7[82],uut.s7[44],uut.s11[20],uut.s11[57],uut.s5[116],uut.s8[15],uut.s5[121],uut.s1[103],uut.s3[101],uut.s10[77],uut.s8[26],uut.s5[119],uut.s7[81],uut.s1[58],uut.s10[70],uut.s1[50],uut.s1[70],uut.s7[80],uut.s11[17],uut.s5[53],uut.s7[126],uut.s1[34],uut.s1[20],uut.s7[56],uut.s6[38],uut.s3[62],uut.s6[102],uut.s9[36],uut.s3[2],uut.s10[75],uut.s1[73],uut.s10[4],uut.s11[64],uut.s2[103],uut.s11[72],uut.s8[76],uut.s3[11],uut.s10[18],uut.s11[63],uut.s5[28],uut.s8[17],uut.s9[44],uut.s5[60],uut.s10[124],uut.s11[31],uut.s3[94],uut.s4[63],uut.s8[73],uut.s9[125],uut.s4[37],uut.s5[114],uut.s3[58],uut.s7[55],uut.s6[72],uut.s5[24],uut.s4[19],uut.s1[92],uut.s3[110],uut.s7[122],uut.s7[106],uut.s8[20],uut.s9[65],uut.s1[13],uut.s10[54],uut.s10[32],uut.s2[104],uut.s3[125],uut.s5[86],uut.s1[65],uut.s6[90],uut.s1[120],uut.s9[20],uut.s9[114],uut.s10[105],uut.s7[124],uut.s9[127],uut.s3[120],uut.s4[86],uut.s10[89],uut.s5[78],uut.s8[118],uut.s2[59],uut.s10[104],uut.s10[58],uut.s6[58],uut.s4[77],uut.s10[85],uut.s6[106],uut.s11[34],uut.s10[29],uut.s11[47],uut.s10[115],uut.s5[37],uut.s11[112],uut.s7[9],uut.s9[75],uut.s11[87],uut.s2[40],uut.s6[83],uut.s2[38],uut.s2[92],uut.s2[106],uut.s9[47],uut.s8[94],uut.s7[31],uut.s1[85],uut.s3[116],uut.s6[65],uut.s2[56],uut.s4[109],uut.s9[26],uut.s10[0],uut.s8[44],uut.s1[127],uut.s5[12],uut.s2[78],uut.s11[124],uut.s8[24],uut.s2[15],uut.s9[78],uut.s11[37],uut.s8[13],uut.s1[1],uut.s11[86],uut.s4[3],uut.s8[72],uut.s11[56],uut.s7[63],uut.s2[21],uut.s3[17],uut.s5[109],uut.s9[2],uut.s3[46],uut.s5[9],uut.s8[50],uut.s3[1],uut.s4[34],uut.s9[32],uut.s8[42],uut.s7[109],uut.s1[37],uut.s1[12],uut.s3[108],uut.s5[99],uut.s5[98],uut.s3[67],uut.s4[59],uut.s5[26],uut.s2[6],uut.s9[8],uut.s10[69],uut.s9[37],uut.s3[93],uut.s10[45],uut.s6[62],uut.s3[77],uut.s1[75],uut.s7[107],uut.s6[108],uut.s8[8],uut.s6[57],uut.s9[58],uut.s1[28],uut.s7[57],uut.s10[109],uut.s7[105],uut.s6[110],uut.s4[30],uut.s6[11],uut.s4[87],uut.s10[56],uut.s6[19],uut.s6[41],uut.s5[38],uut.s8[12],uut.s11[98],uut.s2[29],uut.s2[34],uut.s8[89],uut.s6[14],uut.s2[114],uut.s2[25],uut.s5[64],uut.s11[82],uut.s1[18],uut.s7[43],uut.s9[46],uut.s4[80],uut.s7[108],uut.s11[69],uut.s11[89],uut.s5[39],uut.s9[0],uut.s3[42],uut.s6[42],uut.s6[111],uut.s9[52],uut.s7[26],uut.s1[95],uut.s4[72],uut.s2[41],uut.s2[0],uut.s1[122],uut.s5[35],uut.s6[88],uut.s9[41],uut.s5[40],uut.s4[83],uut.s5[125],uut.s1[77],uut.s8[53],uut.s7[10],uut.s9[64],uut.s6[80],uut.s4[11],uut.s8[107],uut.s10[42],uut.s5[89],uut.s3[6],uut.s6[125],uut.s5[120],uut.s6[74],uut.s2[9],uut.s9[108],uut.s2[26],uut.s3[23],uut.s11[19],uut.s5[82],uut.s6[100],uut.s3[109],uut.s6[7],uut.s10[82],uut.s4[38],uut.s5[110],uut.s3[117],uut.s4[51],uut.s6[0],uut.s9[24],uut.s3[35],uut.s10[111],uut.s2[28],uut.s1[72],uut.s2[48],uut.s2[120],uut.s6[27],uut.s6[73],uut.s8[61],uut.s9[63],uut.s11[40],uut.s8[37],uut.s10[17],uut.s11[29],uut.s7[5],uut.s1[26],uut.s6[86],uut.s5[5],uut.s3[88],uut.s5[106],uut.s7[123],uut.s3[19],uut.s3[57],uut.s1[101],uut.s7[113],uut.s11[92],uut.s7[73],uut.s3[54],uut.s11[74],uut.s11[5],uut.s10[11],uut.s3[45],uut.s3[91],uut.s2[111],uut.s5[44],uut.s4[50],uut.s3[84],uut.s1[40],uut.s2[18],uut.s6[50],uut.s2[49],uut.s7[64],uut.s7[38],uut.s1[100],uut.s4[103],uut.s2[100],uut.s8[92],uut.s11[11],uut.s5[45],uut.s3[119],uut.s1[31],uut.s4[117],uut.s6[112],uut.s2[1],uut.s11[105],uut.s8[2],uut.s4[82],uut.s8[58],uut.s7[120],uut.s9[89],uut.s7[93],uut.s3[114],uut.s9[25],uut.s4[67],uut.s1[59],uut.s7[17],uut.s11[109],uut.s10[24],uut.s1[123],uut.s8[10],uut.s6[117],uut.s11[100],uut.s8[34],uut.s8[104],uut.s8[36],uut.s7[50],uut.s2[79],uut.s1[63],uut.s3[55],uut.s7[104],uut.s6[24],uut.s3[95],uut.s11[14],uut.s8[18],uut.s1[42],uut.s4[13],uut.s1[23],uut.s8[121],uut.s5[88],uut.s8[45],uut.s2[10],uut.s10[113],uut.s6[95],uut.s1[124],uut.s7[86],uut.s1[81],uut.s7[20],uut.s1[17],uut.s11[18],uut.s8[33],uut.s10[118],uut.s8[114],uut.s6[115],uut.s6[66],uut.s4[47],uut.s9[107],uut.s9[21],uut.s11[73],uut.s7[24],uut.s10[8],uut.s3[71],uut.s7[28],uut.s4[41],uut.s7[34],uut.s6[5],uut.s11[96],uut.s8[70],uut.s10[116],uut.s9[119],uut.s8[120],uut.s5[57],uut.s11[115],uut.s9[14],uut.s9[113],uut.s4[81],uut.s11[97],uut.s8[48],uut.s11[0],uut.s4[120],uut.s8[111],uut.s5[63],uut.s10[25],uut.s9[91],uut.s9[121],uut.s11[125],uut.s3[31],uut.s2[53],uut.s11[78],uut.s4[96],uut.s3[102],uut.s6[28],uut.s4[40],uut.s8[43],uut.s2[37],uut.s6[84],uut.s9[86],uut.s4[106],uut.s5[100],uut.s11[62],uut.s4[2],uut.s9[96],uut.s2[95],uut.s4[78],uut.s7[22],uut.s11[39],uut.s5[104],uut.s8[25],uut.s9[56],uut.s10[22],uut.s2[11],uut.s5[62],uut.s5[13],uut.s5[80],uut.s7[99],uut.s10[36],uut.s10[64],uut.s10[14],uut.s7[27],uut.s1[44],uut.s1[114],uut.s7[36],uut.s8[22],uut.s7[2],uut.s1[76],uut.s10[52],uut.s2[39],uut.s10[63],uut.s9[68],uut.s2[57],uut.s4[49],uut.s1[60],uut.s4[23],uut.s11[79],uut.s8[51],uut.s8[100],uut.s5[115],uut.s1[53],uut.s5[1],uut.s1[99],uut.s2[16],uut.s4[21],uut.s4[123],uut.s7[61],uut.s9[100],uut.s1[91],uut.s1[64],uut.s10[80],uut.s10[3],uut.s3[106],uut.s9[74],uut.s10[95],uut.s4[99],uut.s4[127],uut.s8[97],uut.s5[108],uut.s11[68],uut.s7[90],uut.s8[41],uut.s9[101],uut.s4[31],uut.s8[81],uut.s1[98],uut.s11[54],uut.s3[7],uut.s3[72],uut.s10[88],uut.s11[123],uut.s1[71],uut.s5[93],uut.s10[90],uut.s9[61],uut.s3[126],uut.s2[109],uut.s8[46],uut.s6[10],uut.s4[115],uut.s5[3],uut.s2[97],uut.s3[27],uut.s10[83],uut.s9[103],uut.s1[3],uut.s7[77],uut.s10[79],uut.s8[75],uut.s10[10],uut.s5[123],uut.s5[30],uut.s7[13],uut.s8[102],uut.s9[22],uut.s9[82],uut.s5[23],uut.s1[104],uut.s10[120],uut.s8[125],uut.s3[90],uut.s3[70],uut.s10[119],uut.s11[91],uut.s7[114],uut.s4[60],uut.s4[124],uut.s8[101],uut.s6[85],uut.s4[1],uut.s3[48],uut.s4[121],uut.s2[19],uut.s7[39],uut.s7[96],uut.s9[43],uut.s1[94],uut.s11[48],uut.s4[100],uut.s8[4],uut.s7[85],uut.s1[86],uut.s1[78],uut.s2[51],uut.s2[13],uut.s4[20],uut.s7[59],uut.s4[116],uut.s2[115],uut.s5[75],uut.s4[75],uut.s5[41],uut.s2[45],uut.s10[12],uut.s11[102],uut.s4[57],uut.s11[16],uut.s9[71],uut.s2[83],uut.s8[62],uut.s2[102],uut.s2[94],uut.s6[119],uut.s4[119],uut.s6[68],uut.s7[83],uut.s1[47],uut.s11[49],uut.s5[10],uut.s9[54],uut.s11[81],uut.s8[5],uut.s4[16],uut.s5[91],uut.s9[51],uut.s6[63],uut.s3[76],uut.s1[96],uut.s5[66],uut.s7[46],uut.s10[2],uut.s7[115],uut.s2[42],uut.s8[112],uut.s10[37],uut.s2[20],uut.s2[35],uut.s11[6],uut.s7[51],uut.s3[38],uut.s11[28],uut.s4[52],uut.s1[107],uut.s4[24],uut.s8[106],uut.s8[28],uut.s6[70],uut.s8[56],uut.s9[5],uut.s4[32],uut.s6[12],uut.s8[40],uut.s2[4],uut.s9[123],uut.s8[9],uut.s10[126],uut.s1[49],uut.s7[12],uut.s11[116],uut.s6[116],uut.s3[40],uut.s5[67],uut.s6[118],uut.s8[105],uut.s1[5],uut.s5[118],uut.s9[31],uut.s3[22],uut.s3[78],uut.s11[118],uut.s3[52],uut.s4[22],uut.s1[14],uut.s8[74],uut.s9[1],uut.s5[51],uut.s9[17],uut.s4[27],uut.s1[115],uut.s9[90],uut.s3[4],uut.s4[48],uut.s9[6],uut.s6[44],uut.s6[20],uut.s5[52],uut.s2[7],uut.s8[39],uut.s3[51],uut.s10[117],uut.s7[48],uut.s4[18],uut.s8[123],uut.s9[23],uut.s6[96],uut.s7[87],uut.s8[57],uut.s2[105],uut.s2[68],uut.s2[80],uut.s2[3],uut.s5[74],uut.s3[44],uut.s4[46],uut.s3[24],uut.s11[7],uut.s3[60],uut.s1[116],uut.s7[103],uut.s9[83],uut.s8[99],uut.s10[60],uut.s10[101],uut.s5[112],uut.s7[110],uut.s6[35],uut.s3[80],uut.s6[123],uut.s10[72],uut.s2[110],uut.s8[64],uut.s11[101],uut.s9[3],uut.s6[77],uut.s10[121],uut.s10[55],uut.s5[17],uut.s2[5],uut.s3[69],uut.s9[28],uut.s4[26],uut.s7[4],uut.s8[116],uut.s7[35],uut.s9[120],uut.s6[6],uut.s5[49],uut.s4[114],uut.s4[17],uut.s11[71],uut.s2[81],uut.s3[41],uut.s6[22],uut.s7[95],uut.s5[81],uut.s8[119],uut.s6[121],uut.s3[112],uut.s11[4],uut.s6[43],uut.s9[126],uut.s10[81],uut.s6[82],uut.s3[63],uut.s6[93],uut.s6[89],uut.s1[68],uut.s7[102],uut.s1[2],uut.s5[90],uut.s6[23],uut.s5[46],uut.s9[60],uut.s11[114],uut.s1[30],uut.s3[107],uut.s4[15],uut.s3[122],uut.s1[36],uut.s4[45],uut.s3[8],uut.s5[0],uut.s6[52],uut.s3[0],uut.s4[71],uut.s2[36],uut.s5[71],uut.s4[122],uut.s1[112],uut.s5[79],uut.s9[19],uut.s3[43],uut.s10[20],uut.s7[119],uut.s1[121],uut.s2[23],uut.s7[1],uut.s7[11],uut.s9[42],uut.s11[36],uut.s4[36],uut.s2[113],uut.s4[126],uut.s9[106],uut.s7[33],uut.s11[45],uut.s5[59],uut.s5[102],uut.s3[73],uut.s11[95],uut.s2[2],uut.s11[110],uut.s6[16],uut.s3[85],uut.s10[114],uut.s5[6],uut.s3[104],uut.s9[9],uut.s10[41],uut.s2[117],uut.s7[29],uut.s1[22],uut.s2[108],uut.s5[54],uut.s6[104],uut.s3[30],uut.s1[24],uut.s7[45],uut.s8[29],uut.s11[26],uut.s2[17],uut.s7[118],uut.s6[34],uut.s5[72],uut.s6[26],uut.s9[79],uut.s6[60],uut.s2[66],uut.s5[101],uut.s4[12],uut.s4[104],uut.s11[51],uut.s4[110],uut.s4[74],uut.s6[91],uut.s8[93],uut.s10[53],uut.s7[84],uut.s4[79],uut.s4[56],uut.s10[67],uut.s7[117],uut.s3[118],uut.s9[66],uut.s11[53],uut.s5[105],uut.s2[50],uut.s5[69],uut.s3[87],uut.s9[16],uut.s8[65],uut.s7[54],uut.s10[97],uut.s3[115],uut.s9[39],uut.s6[8],uut.s8[63],uut.s8[27],uut.s8[30],uut.s3[14],uut.s5[15],uut.s10[122],uut.s10[23],uut.s5[95],uut.s9[92],uut.s7[14],uut.s11[10],uut.s1[61],uut.s5[16],uut.s1[4],uut.s10[46],uut.s1[84],uut.s9[102],uut.s10[108],uut.s7[74],uut.s9[48],uut.s2[99],uut.s4[44],uut.s3[47],uut.s11[84],uut.s10[73],uut.s7[65],uut.s7[75],uut.s1[88],uut.s6[21],uut.s2[32],uut.s4[90],uut.s8[69],uut.s5[77],uut.s1[118],uut.s2[86],uut.s3[66],uut.s1[113],uut.s10[48],uut.s4[8],uut.s5[11],uut.s3[33],uut.s6[87],uut.s6[9],uut.s5[97],uut.s9[122],uut.s10[50],uut.s9[45],uut.s6[79],uut.s2[84],uut.s1[27],uut.s10[66],uut.s1[74],uut.s7[15],uut.s2[107],uut.s4[105],uut.s5[76],uut.s9[59],uut.s4[91],uut.s6[3],uut.s8[108],uut.s3[37],uut.s11[52],uut.s2[60],uut.s7[49],uut.s7[41],uut.s6[25],uut.s6[29],uut.s10[43],uut.s4[35],uut.s7[71],uut.s8[95],uut.s5[22],uut.s1[69],uut.s6[54],uut.s3[49],uut.s5[50],uut.s2[73],uut.s6[32],uut.s2[118],uut.s11[65],uut.s2[12],uut.s6[127],uut.s5[32],uut.s1[51],uut.s2[67],uut.s9[94],uut.s9[53],uut.s9[118],uut.s9[97],uut.s1[80],uut.s5[85],uut.s6[69],uut.s5[4],uut.s9[50],uut.s11[35],uut.s11[88],uut.s11[59],uut.s1[105],uut.s8[86],uut.s1[57],uut.s6[40],uut.s1[10],uut.s1[29],uut.s8[55],uut.s8[52],uut.s5[113],uut.s10[84],uut.s11[9],uut.s2[125],uut.s9[10],uut.s1[19],uut.s5[27],uut.s7[121],uut.s11[99],uut.s5[58],uut.s5[8],uut.s8[23],uut.s11[50],uut.s10[76],uut.s3[81],uut.s2[116],uut.s3[13],uut.s7[32],uut.s9[12],uut.s3[68],uut.s11[43],uut.s1[89],uut.s7[94],uut.s2[112],uut.s3[64],uut.s4[39],uut.s5[14],uut.s6[31],uut.s7[116],uut.s4[102],uut.s4[84],uut.s2[76],uut.s9[7],uut.s10[49],uut.s10[106],uut.s9[111],uut.s10[125],uut.s10[65],uut.s5[33],uut.s11[46],uut.s2[82],uut.s9[95],uut.s6[13],uut.s10[51],uut.s6[17],uut.s1[21],uut.s2[93],uut.s2[14],uut.s7[88],uut.s9[72],uut.s11[117],uut.s11[94],uut.s8[38],uut.s4[94],uut.s6[99],uut.s6[47],uut.s11[127],uut.s2[119],uut.s5[56],uut.s1[79],uut.s10[92],uut.s4[64],uut.s1[7],uut.s7[3],uut.s11[55],uut.s4[33],uut.s2[124],uut.s7[53],uut.s9[38],uut.s10[78],uut.s11[12],uut.s10[9],uut.s7[100],uut.s4[42],uut.s2[47],uut.s10[91],uut.s10[103],uut.s10[33],uut.s8[98],uut.s1[9],uut.s8[59],uut.s11[27],uut.s3[100],uut.s3[79],uut.s8[77],uut.s3[98],uut.s8[11],uut.s3[5],uut.s4[9],uut.s9[33],uut.s11[66],uut.s11[76],uut.s2[75],uut.s4[68],uut.s10[107],uut.s6[30],uut.s11[3],uut.s5[96],uut.s7[97],uut.s11[2],uut.s8[14],uut.s5[126],uut.s3[89],uut.s6[39],uut.s4[89],uut.s6[64],uut.s8[80],uut.s1[125],uut.s4[66],uut.s11[25],uut.s4[62],uut.s8[84],uut.s3[61],uut.s4[93],uut.s7[69],uut.s9[27],uut.s4[5],uut.s4[28],uut.s10[87],uut.s1[126],uut.s4[98],uut.s7[91],uut.s6[113],uut.s7[21],uut.s9[117],uut.s5[31],uut.s2[22],uut.s5[47],uut.s5[55],uut.s4[97],uut.s11[113],uut.s8[113],uut.s6[124],uut.s9[73],uut.s3[29],uut.s5[103],uut.s8[7],uut.s8[115],uut.s10[19],uut.s4[29],uut.s2[89],uut.s10[15],uut.s2[55],uut.s4[6],uut.s11[13],uut.s11[80],uut.s3[39],uut.s10[102],uut.s1[102],uut.s2[46],uut.s4[58],uut.s6[49],uut.s8[60],uut.s10[35],uut.s7[62],uut.s11[122],uut.s1[109],uut.s3[28],uut.s8[68],uut.s10[31],uut.s10[57],uut.s8[35],uut.s3[32],uut.s9[80],uut.s8[3],uut.s8[49],uut.s2[54],uut.s6[97],uut.s4[108],uut.s11[111],uut.s10[62],uut.s10[61],uut.s10[5],uut.s2[77],uut.s5[2],uut.s4[73],uut.s5[36],uut.s7[127],uut.s2[127],uut.s8[110],uut.s10[112],uut.s11[22],uut.s7[8],uut.s6[37],uut.s2[91],uut.s7[112],uut.s5[42],uut.s4[88],uut.s8[122],uut.s2[65],uut.s9[77],uut.s8[47],uut.s11[119],uut.s3[65],uut.s2[58],uut.s6[107],uut.s6[56],uut.s10[39],uut.s2[74],uut.s3[97],uut.s10[30],uut.s9[124],uut.s7[23],uut.s11[120],uut.s6[59],uut.s1[119],uut.s9[18],uut.s7[79],uut.s2[123],uut.s6[120],uut.s3[105],uut.s3[36],uut.s3[99],uut.s2[69],uut.s8[82],uut.s2[64],uut.s3[103],uut.s1[67],uut.s1[35],uut.s7[76],uut.s5[84],uut.s10[16],uut.s9[109],uut.s11[60],uut.s6[92],uut.s2[8],uut.s7[0],uut.s5[18],uut.s5[21],uut.s10[68],uut.s7[70],uut.s5[124],uut.s10[98],uut.s3[111],uut.s1[48],uut.s9[70],uut.s7[7],uut.s6[4],uut.s1[0],uut.s10[93],uut.s6[51],uut.s10[26],uut.s7[111],uut.s2[85],uut.s4[65],uut.s3[92],uut.s9[99],uut.s6[36],uut.s8[117],uut.s7[16],uut.s10[6],uut.s8[16],uut.s4[25],uut.s6[98],uut.s2[101],uut.s11[103],uut.s11[23],uut.s11[8],uut.s5[48],uut.s1[6],uut.s1[110],uut.s10[59],uut.s8[66],uut.s11[15],uut.s1[8],uut.s10[27],uut.s2[61],uut.s5[111],uut.s6[71],uut.s10[94],uut.s11[21],uut.s11[30],uut.s7[19],uut.s10[7],uut.s11[67],uut.s4[54],uut.s7[125],uut.s1[97],uut.s11[58],uut.s6[2],uut.s11[38],uut.s4[85],uut.s8[85],uut.s10[74],uut.s8[126],uut.s4[55],uut.s7[18],uut.s8[103],uut.s4[95],uut.s3[20],uut.s1[46],uut.s10[127],uut.s1[16],uut.s5[65],uut.s8[127],uut.s7[40],uut.s3[83],uut.s9[85],uut.s4[14],uut.s2[30],uut.s11[93],uut.s3[34],uut.s5[83],uut.s9[30],uut.s8[87],uut.s3[121],uut.s4[0],uut.s1[117],uut.s7[42],uut.s11[85],uut.s5[127],uut.s4[70],uut.s6[53],uut.s2[121],uut.s4[76],uut.s6[67],uut.s3[50],uut.s1[83],uut.s10[13],uut.s7[58],uut.s10[34],uut.s7[37],uut.s6[114],uut.s4[7],uut.s10[99],uut.s4[4],uut.s8[79],uut.s3[74],uut.s9[35],uut.s9[15],uut.s11[1],uut.s3[124],uut.s2[72],uut.s1[32],uut.s9[105],uut.s10[1],uut.s9[84],uut.s11[121],uut.s6[15],uut.s6[61],uut.s3[21],uut.s1[93],uut.s5[20],uut.s9[29],uut.s5[29],uut.s2[63],uut.s9[4],uut.s8[90],uut.s1[55],uut.s1[11],uut.s3[15],uut.s6[126],uut.s1[87],uut.s3[12],uut.s5[94],uut.s7[92],uut.s7[72],uut.s8[31],uut.s11[24],uut.s2[87],uut.s2[98],uut.s3[3],uut.s6[48],uut.s7[98],uut.s4[92],uut.s2[44],uut.s1[25],uut.s11[61],uut.s7[6],uut.s5[73],uut.s7[30],uut.s10[71],uut.s6[81],uut.s1[45],uut.s2[122],uut.s9[112],uut.s6[103],uut.s6[76],uut.s9[93],uut.s10[123],uut.s3[56],uut.s11[41],uut.s11[42],uut.s3[127],uut.s3[26],uut.s10[86],uut.s10[47],uut.s1[66],uut.s5[7],uut.s5[70],uut.s3[123],uut.s10[110],uut.s11[83],uut.s3[53],uut.s6[45],uut.s2[71],uut.s9[11],uut.s1[106],uut.s6[33],uut.s5[107],uut.s4[10],uut.s3[113]};
			//data1 <= data1_1;

		end


		always@(posedge clk)
		begin
			if(rst)
    data2<= 0;
			else
    data2<=data1;
	 //data2 <= data2_1;
		end		

		
		reg signed [15:0]plot;
		always@(posedge clk)
		begin
			if(rst)
    plot<= 0;
		else
		plot<= (64*(data2[1407]^data1[1407])+2*(data2[1406]^data1[1406])+64*(data2[1405]^data1[1405])+64*(data2[1404]^data1[1404])+16*(data2[1403]^data1[1403])+64*(data2[1402]^data1[1402])+64*(data2[1401]^data1[1401])+2*(data2[1400]^data1[1400])+2*(data2[1399]^data1[1399])+64*(data2[1398]^data1[1398])+16*(data2[1397]^data1[1397])+32*(data2[1396]^data1[1396])+32*(data2[1395]^data1[1395])+2*(data2[1394]^data1[1394])+2*(data2[1393]^data1[1393])+2*(data2[1392]^data1[1392])+64*(data2[1391]^data1[1391])+64*(data2[1390]^data1[1390])+33*(data2[1389]^data1[1389])+2*(data2[1388]^data1[1388])+2*(data2[1387]^data1[1387])+32*(data2[1386]^data1[1386])+2*(data2[1385]^data1[1385])+64*(data2[1384]^data1[1384])+32*(data2[1383]^data1[1383])+2*(data2[1382]^data1[1382])+64*(data2[1381]^data1[1381])+64*(data2[1380]^data1[1380])+2*(data2[1379]^data1[1379])+2*(data2[1378]^data1[1378])+2*(data2[1377]^data1[1377])+2*(data2[1376]^data1[1376])+2*(data2[1375]^data1[1375])+33*(data2[1374]^data1[1374])+2*(data2[1373]^data1[1373])+64*(data2[1372]^data1[1372])+32*(data2[1371]^data1[1371])+64*(data2[1370]^data1[1370])+64*(data2[1369]^data1[1369])+2*(data2[1368]^data1[1368])+16*(data2[1367]^data1[1367])+64*(data2[1366]^data1[1366])+2*(data2[1365]^data1[1365])+64*(data2[1364]^data1[1364])+64*(data2[1363]^data1[1363])+2*(data2[1362]^data1[1362])+2*(data2[1361]^data1[1361])+33*(data2[1360]^data1[1360])+2*(data2[1359]^data1[1359])+2*(data2[1358]^data1[1358])+9*(data2[1357]^data1[1357])+33*(data2[1356]^data1[1356])+2*(data2[1355]^data1[1355])+2*(data2[1354]^data1[1354])+33*(data2[1353]^data1[1353])+32*(data2[1352]^data1[1352])+32*(data2[1351]^data1[1351])+64*(data2[1350]^data1[1350])+32*(data2[1349]^data1[1349])+64*(data2[1348]^data1[1348])+2*(data2[1347]^data1[1347])+64*(data2[1346]^data1[1346])+2*(data2[1345]^data1[1345])+2*(data2[1344]^data1[1344])+64*(data2[1343]^data1[1343])+64*(data2[1342]^data1[1342])+2*(data2[1341]^data1[1341])+33*(data2[1340]^data1[1340])+2*(data2[1339]^data1[1339])+32*(data2[1338]^data1[1338])+64*(data2[1337]^data1[1337])+64*(data2[1336]^data1[1336])+2*(data2[1335]^data1[1335])+2*(data2[1334]^data1[1334])+16*(data2[1333]^data1[1333])+64*(data2[1332]^data1[1332])+2*(data2[1331]^data1[1331])+2*(data2[1330]^data1[1330])+2*(data2[1329]^data1[1329])+2*(data2[1328]^data1[1328])+2*(data2[1327]^data1[1327])+32*(data2[1326]^data1[1326])+2*(data2[1325]^data1[1325])+64*(data2[1324]^data1[1324])+32*(data2[1323]^data1[1323])+2*(data2[1322]^data1[1322])+2*(data2[1321]^data1[1321])+2*(data2[1320]^data1[1320])+32*(data2[1319]^data1[1319])+64*(data2[1318]^data1[1318])+2*(data2[1317]^data1[1317])+32*(data2[1316]^data1[1316])+2*(data2[1315]^data1[1315])+2*(data2[1314]^data1[1314])+32*(data2[1313]^data1[1313])+2*(data2[1312]^data1[1312])+64*(data2[1311]^data1[1311])+2*(data2[1310]^data1[1310])+32*(data2[1309]^data1[1309])+64*(data2[1308]^data1[1308])+32*(data2[1307]^data1[1307])+2*(data2[1306]^data1[1306])+2*(data2[1305]^data1[1305])+16*(data2[1304]^data1[1304])+64*(data2[1303]^data1[1303])+64*(data2[1302]^data1[1302])+33*(data2[1301]^data1[1301])+2*(data2[1300]^data1[1300])+64*(data2[1299]^data1[1299])+64*(data2[1298]^data1[1298])+2*(data2[1297]^data1[1297])+2*(data2[1296]^data1[1296])+2*(data2[1295]^data1[1295])+64*(data2[1294]^data1[1294])+32*(data2[1293]^data1[1293])+2*(data2[1292]^data1[1292])+2*(data2[1291]^data1[1291])+2*(data2[1290]^data1[1290])+2*(data2[1289]^data1[1289])+2*(data2[1288]^data1[1288])+16*(data2[1287]^data1[1287])+16*(data2[1286]^data1[1286])+2*(data2[1285]^data1[1285])+2*(data2[1284]^data1[1284])+2*(data2[1283]^data1[1283])+2*(data2[1282]^data1[1282])+2*(data2[1281]^data1[1281])+32*(data2[1280]^data1[1280])+64*(data2[1279]^data1[1279])+64*(data2[1278]^data1[1278])+2*(data2[1277]^data1[1277])+2*(data2[1276]^data1[1276])+2*(data2[1275]^data1[1275])+32*(data2[1274]^data1[1274])+32*(data2[1273]^data1[1273])+33*(data2[1272]^data1[1272])+2*(data2[1271]^data1[1271])+33*(data2[1270]^data1[1270])+64*(data2[1269]^data1[1269])+64*(data2[1268]^data1[1268])+2*(data2[1267]^data1[1267])+2*(data2[1266]^data1[1266])+9*(data2[1265]^data1[1265])+2*(data2[1264]^data1[1264])+64*(data2[1263]^data1[1263])+2*(data2[1262]^data1[1262])+64*(data2[1261]^data1[1261])+32*(data2[1260]^data1[1260])+2*(data2[1259]^data1[1259])+32*(data2[1258]^data1[1258])+33*(data2[1257]^data1[1257])+2*(data2[1256]^data1[1256])+64*(data2[1255]^data1[1255])+64*(data2[1254]^data1[1254])+2*(data2[1253]^data1[1253])+2*(data2[1252]^data1[1252])+32*(data2[1251]^data1[1251])+2*(data2[1250]^data1[1250])+2*(data2[1249]^data1[1249])+64*(data2[1248]^data1[1248])+2*(data2[1247]^data1[1247])+64*(data2[1246]^data1[1246])+2*(data2[1245]^data1[1245])+32*(data2[1244]^data1[1244])+64*(data2[1243]^data1[1243])+32*(data2[1242]^data1[1242])+2*(data2[1241]^data1[1241])+64*(data2[1240]^data1[1240])+2*(data2[1239]^data1[1239])+8*(data2[1238]^data1[1238])+64*(data2[1237]^data1[1237])+2*(data2[1236]^data1[1236])+2*(data2[1235]^data1[1235])+33*(data2[1234]^data1[1234])+2*(data2[1233]^data1[1233])+8*(data2[1232]^data1[1232])+32*(data2[1231]^data1[1231])+16*(data2[1230]^data1[1230])+2*(data2[1229]^data1[1229])+2*(data2[1228]^data1[1228])+64*(data2[1227]^data1[1227])+33*(data2[1226]^data1[1226])+64*(data2[1225]^data1[1225])+2*(data2[1224]^data1[1224])+2*(data2[1223]^data1[1223])+64*(data2[1222]^data1[1222])+64*(data2[1221]^data1[1221])+64*(data2[1220]^data1[1220])+32*(data2[1219]^data1[1219])+2*(data2[1218]^data1[1218])+2*(data2[1217]^data1[1217])+2*(data2[1216]^data1[1216])+2*(data2[1215]^data1[1215])+64*(data2[1214]^data1[1214])+2*(data2[1213]^data1[1213])+2*(data2[1212]^data1[1212])+64*(data2[1211]^data1[1211])+64*(data2[1210]^data1[1210])+17*(data2[1209]^data1[1209])+64*(data2[1208]^data1[1208])+2*(data2[1207]^data1[1207])+64*(data2[1206]^data1[1206])+2*(data2[1205]^data1[1205])+2*(data2[1204]^data1[1204])+2*(data2[1203]^data1[1203])+2*(data2[1202]^data1[1202])+2*(data2[1201]^data1[1201])+64*(data2[1200]^data1[1200])+32*(data2[1199]^data1[1199])+2*(data2[1198]^data1[1198])+17*(data2[1197]^data1[1197])+2*(data2[1196]^data1[1196])+64*(data2[1195]^data1[1195])+2*(data2[1194]^data1[1194])+2*(data2[1193]^data1[1193])+2*(data2[1192]^data1[1192])+64*(data2[1191]^data1[1191])+2*(data2[1190]^data1[1190])+2*(data2[1189]^data1[1189])+32*(data2[1188]^data1[1188])+2*(data2[1187]^data1[1187])+8*(data2[1186]^data1[1186])+2*(data2[1185]^data1[1185])+33*(data2[1184]^data1[1184])+32*(data2[1183]^data1[1183])+2*(data2[1182]^data1[1182])+2*(data2[1181]^data1[1181])+8*(data2[1180]^data1[1180])+64*(data2[1179]^data1[1179])+2*(data2[1178]^data1[1178])+32*(data2[1177]^data1[1177])+64*(data2[1176]^data1[1176])+64*(data2[1175]^data1[1175])+2*(data2[1174]^data1[1174])+2*(data2[1173]^data1[1173])+2*(data2[1172]^data1[1172])+64*(data2[1171]^data1[1171])+64*(data2[1170]^data1[1170])+2*(data2[1169]^data1[1169])+64*(data2[1168]^data1[1168])+64*(data2[1167]^data1[1167])+2*(data2[1166]^data1[1166])+2*(data2[1165]^data1[1165])+2*(data2[1164]^data1[1164])+16*(data2[1163]^data1[1163])+64*(data2[1162]^data1[1162])+32*(data2[1161]^data1[1161])+32*(data2[1160]^data1[1160])+2*(data2[1159]^data1[1159])+64*(data2[1158]^data1[1158])+2*(data2[1157]^data1[1157])+32*(data2[1156]^data1[1156])+2*(data2[1155]^data1[1155])+64*(data2[1154]^data1[1154])+16*(data2[1153]^data1[1153])+64*(data2[1152]^data1[1152])+2*(data2[1151]^data1[1151])+32*(data2[1150]^data1[1150])+2*(data2[1149]^data1[1149])+64*(data2[1148]^data1[1148])+64*(data2[1147]^data1[1147])+33*(data2[1146]^data1[1146])+2*(data2[1145]^data1[1145])+32*(data2[1144]^data1[1144])+16*(data2[1143]^data1[1143])+2*(data2[1142]^data1[1142])+64*(data2[1141]^data1[1141])+64*(data2[1140]^data1[1140])+2*(data2[1139]^data1[1139])+2*(data2[1138]^data1[1138])+2*(data2[1137]^data1[1137])+64*(data2[1136]^data1[1136])+64*(data2[1135]^data1[1135])+64*(data2[1134]^data1[1134])+9*(data2[1133]^data1[1133])+17*(data2[1132]^data1[1132])+64*(data2[1131]^data1[1131])+64*(data2[1130]^data1[1130])+64*(data2[1129]^data1[1129])+32*(data2[1128]^data1[1128])+2*(data2[1127]^data1[1127])+2*(data2[1126]^data1[1126])+2*(data2[1125]^data1[1125])+64*(data2[1124]^data1[1124])+2*(data2[1123]^data1[1123])+2*(data2[1122]^data1[1122])+64*(data2[1121]^data1[1121])+64*(data2[1120]^data1[1120])+2*(data2[1119]^data1[1119])+2*(data2[1118]^data1[1118])+2*(data2[1117]^data1[1117])+2*(data2[1116]^data1[1116])+2*(data2[1115]^data1[1115])+64*(data2[1114]^data1[1114])+2*(data2[1113]^data1[1113])+2*(data2[1112]^data1[1112])+2*(data2[1111]^data1[1111])+2*(data2[1110]^data1[1110])+32*(data2[1109]^data1[1109])+2*(data2[1108]^data1[1108])+16*(data2[1107]^data1[1107])+2*(data2[1106]^data1[1106])+2*(data2[1105]^data1[1105])+2*(data2[1104]^data1[1104])+17*(data2[1103]^data1[1103])+2*(data2[1102]^data1[1102])+16*(data2[1101]^data1[1101])+64*(data2[1100]^data1[1100])+64*(data2[1099]^data1[1099])+2*(data2[1098]^data1[1098])+2*(data2[1097]^data1[1097])+64*(data2[1096]^data1[1096])+64*(data2[1095]^data1[1095])+33*(data2[1094]^data1[1094])+32*(data2[1093]^data1[1093])+64*(data2[1092]^data1[1092])+2*(data2[1091]^data1[1091])+2*(data2[1090]^data1[1090])+64*(data2[1089]^data1[1089])+2*(data2[1088]^data1[1088])+32*(data2[1087]^data1[1087])+32*(data2[1086]^data1[1086])+9*(data2[1085]^data1[1085])+2*(data2[1084]^data1[1084])+64*(data2[1083]^data1[1083])+2*(data2[1082]^data1[1082])+2*(data2[1081]^data1[1081])+2*(data2[1080]^data1[1080])+2*(data2[1079]^data1[1079])+16*(data2[1078]^data1[1078])+64*(data2[1077]^data1[1077])+64*(data2[1076]^data1[1076])+64*(data2[1075]^data1[1075])+64*(data2[1074]^data1[1074])+33*(data2[1073]^data1[1073])+2*(data2[1072]^data1[1072])+2*(data2[1071]^data1[1071])+33*(data2[1070]^data1[1070])+64*(data2[1069]^data1[1069])+33*(data2[1068]^data1[1068])+64*(data2[1067]^data1[1067])+2*(data2[1066]^data1[1066])+2*(data2[1065]^data1[1065])+2*(data2[1064]^data1[1064])+2*(data2[1063]^data1[1063])+64*(data2[1062]^data1[1062])+2*(data2[1061]^data1[1061])+2*(data2[1060]^data1[1060])+33*(data2[1059]^data1[1059])+32*(data2[1058]^data1[1058])+2*(data2[1057]^data1[1057])+33*(data2[1056]^data1[1056])+2*(data2[1055]^data1[1055])+16*(data2[1054]^data1[1054])+2*(data2[1053]^data1[1053])+64*(data2[1052]^data1[1052])+16*(data2[1051]^data1[1051])+32*(data2[1050]^data1[1050])+33*(data2[1049]^data1[1049])+2*(data2[1048]^data1[1048])+64*(data2[1047]^data1[1047])+2*(data2[1046]^data1[1046])+2*(data2[1045]^data1[1045])+32*(data2[1044]^data1[1044])+17*(data2[1043]^data1[1043])+64*(data2[1042]^data1[1042])+64*(data2[1041]^data1[1041])+2*(data2[1040]^data1[1040])+2*(data2[1039]^data1[1039])+64*(data2[1038]^data1[1038])+2*(data2[1037]^data1[1037])+64*(data2[1036]^data1[1036])+64*(data2[1035]^data1[1035])+64*(data2[1034]^data1[1034])+64*(data2[1033]^data1[1033])+2*(data2[1032]^data1[1032])+2*(data2[1031]^data1[1031])+2*(data2[1030]^data1[1030])+2*(data2[1029]^data1[1029])+32*(data2[1028]^data1[1028])+2*(data2[1027]^data1[1027])+2*(data2[1026]^data1[1026])+32*(data2[1025]^data1[1025])+2*(data2[1024]^data1[1024])+64*(data2[1023]^data1[1023])+2*(data2[1022]^data1[1022])+64*(data2[1021]^data1[1021])+64*(data2[1020]^data1[1020])+33*(data2[1019]^data1[1019])+2*(data2[1018]^data1[1018])+64*(data2[1017]^data1[1017])+64*(data2[1016]^data1[1016])+64*(data2[1015]^data1[1015])+2*(data2[1014]^data1[1014])+32*(data2[1013]^data1[1013])+2*(data2[1012]^data1[1012])+32*(data2[1011]^data1[1011])+32*(data2[1010]^data1[1010])+32*(data2[1009]^data1[1009])+2*(data2[1008]^data1[1008])+64*(data2[1007]^data1[1007])+64*(data2[1006]^data1[1006])+16*(data2[1005]^data1[1005])+33*(data2[1004]^data1[1004])+64*(data2[1003]^data1[1003])+64*(data2[1002]^data1[1002])+64*(data2[1001]^data1[1001])+64*(data2[1000]^data1[1000])+2*(data2[999]^data1[999])+64*(data2[998]^data1[998])+2*(data2[997]^data1[997])+2*(data2[996]^data1[996])+64*(data2[995]^data1[995])+64*(data2[994]^data1[994])+64*(data2[993]^data1[993])+2*(data2[992]^data1[992])+32*(data2[991]^data1[991])+33*(data2[990]^data1[990])+16*(data2[989]^data1[989])+16*(data2[988]^data1[988])+64*(data2[987]^data1[987])+2*(data2[986]^data1[986])+64*(data2[985]^data1[985])+32*(data2[984]^data1[984])+2*(data2[983]^data1[983])+64*(data2[982]^data1[982])+2*(data2[981]^data1[981])+2*(data2[980]^data1[980])+2*(data2[979]^data1[979])+2*(data2[978]^data1[978])+64*(data2[977]^data1[977])+2*(data2[976]^data1[976])+64*(data2[975]^data1[975])+64*(data2[974]^data1[974])+2*(data2[973]^data1[973])+32*(data2[972]^data1[972])+2*(data2[971]^data1[971])+64*(data2[970]^data1[970])+2*(data2[969]^data1[969])+2*(data2[968]^data1[968])+32*(data2[967]^data1[967])+2*(data2[966]^data1[966])+2*(data2[965]^data1[965])+2*(data2[964]^data1[964])+2*(data2[963]^data1[963])+16*(data2[962]^data1[962])+16*(data2[961]^data1[961])+16*(data2[960]^data1[960])+2*(data2[959]^data1[959])+2*(data2[958]^data1[958])+16*(data2[957]^data1[957])+32*(data2[956]^data1[956])+2*(data2[955]^data1[955])+64*(data2[954]^data1[954])+64*(data2[953]^data1[953])+16*(data2[952]^data1[952])+2*(data2[951]^data1[951])+33*(data2[950]^data1[950])+2*(data2[949]^data1[949])+64*(data2[948]^data1[948])+2*(data2[947]^data1[947])+2*(data2[946]^data1[946])+64*(data2[945]^data1[945])+2*(data2[944]^data1[944])+64*(data2[943]^data1[943])+2*(data2[942]^data1[942])+64*(data2[941]^data1[941])+32*(data2[940]^data1[940])+2*(data2[939]^data1[939])+2*(data2[938]^data1[938])+2*(data2[937]^data1[937])+2*(data2[936]^data1[936])+2*(data2[935]^data1[935])+16*(data2[934]^data1[934])+2*(data2[933]^data1[933])+2*(data2[932]^data1[932])+32*(data2[931]^data1[931])+2*(data2[930]^data1[930])+2*(data2[929]^data1[929])+16*(data2[928]^data1[928])+2*(data2[927]^data1[927])+64*(data2[926]^data1[926])+2*(data2[925]^data1[925])+2*(data2[924]^data1[924])+32*(data2[923]^data1[923])+2*(data2[922]^data1[922])+2*(data2[921]^data1[921])+2*(data2[920]^data1[920])+2*(data2[919]^data1[919])+33*(data2[918]^data1[918])+32*(data2[917]^data1[917])+2*(data2[916]^data1[916])+2*(data2[915]^data1[915])+64*(data2[914]^data1[914])+32*(data2[913]^data1[913])+2*(data2[912]^data1[912])+32*(data2[911]^data1[911])+64*(data2[910]^data1[910])+2*(data2[909]^data1[909])+9*(data2[908]^data1[908])+2*(data2[907]^data1[907])+2*(data2[906]^data1[906])+2*(data2[905]^data1[905])+32*(data2[904]^data1[904])+16*(data2[903]^data1[903])+64*(data2[902]^data1[902])+16*(data2[901]^data1[901])+64*(data2[900]^data1[900])+64*(data2[899]^data1[899])+2*(data2[898]^data1[898])+64*(data2[897]^data1[897])+2*(data2[896]^data1[896])+64*(data2[895]^data1[895])+2*(data2[894]^data1[894])+2*(data2[893]^data1[893])+64*(data2[892]^data1[892])+33*(data2[891]^data1[891])+16*(data2[890]^data1[890])+64*(data2[889]^data1[889])+2*(data2[888]^data1[888])+16*(data2[887]^data1[887])+32*(data2[886]^data1[886])+2*(data2[885]^data1[885])+8*(data2[884]^data1[884])+33*(data2[883]^data1[883])+2*(data2[882]^data1[882])+2*(data2[881]^data1[881])+2*(data2[880]^data1[880])+64*(data2[879]^data1[879])+17*(data2[878]^data1[878])+64*(data2[877]^data1[877])+33*(data2[876]^data1[876])+2*(data2[875]^data1[875])+2*(data2[874]^data1[874])+2*(data2[873]^data1[873])+2*(data2[872]^data1[872])+2*(data2[871]^data1[871])+64*(data2[870]^data1[870])+64*(data2[869]^data1[869])+2*(data2[868]^data1[868])+2*(data2[867]^data1[867])+2*(data2[866]^data1[866])+64*(data2[865]^data1[865])+2*(data2[864]^data1[864])+16*(data2[863]^data1[863])+2*(data2[862]^data1[862])+2*(data2[861]^data1[861])+64*(data2[860]^data1[860])+64*(data2[859]^data1[859])+64*(data2[858]^data1[858])+16*(data2[857]^data1[857])+8*(data2[856]^data1[856])+2*(data2[855]^data1[855])+2*(data2[854]^data1[854])+33*(data2[853]^data1[853])+64*(data2[852]^data1[852])+64*(data2[851]^data1[851])+16*(data2[850]^data1[850])+64*(data2[849]^data1[849])+64*(data2[848]^data1[848])+64*(data2[847]^data1[847])+2*(data2[846]^data1[846])+2*(data2[845]^data1[845])+64*(data2[844]^data1[844])+64*(data2[843]^data1[843])+2*(data2[842]^data1[842])+2*(data2[841]^data1[841])+64*(data2[840]^data1[840])+2*(data2[839]^data1[839])+2*(data2[838]^data1[838])+16*(data2[837]^data1[837])+16*(data2[836]^data1[836])+2*(data2[835]^data1[835])+33*(data2[834]^data1[834])+32*(data2[833]^data1[833])+2*(data2[832]^data1[832])+2*(data2[831]^data1[831])+2*(data2[830]^data1[830])+16*(data2[829]^data1[829])+2*(data2[828]^data1[828])+32*(data2[827]^data1[827])+16*(data2[826]^data1[826])+16*(data2[825]^data1[825])+64*(data2[824]^data1[824])+2*(data2[823]^data1[823])+32*(data2[822]^data1[822])+16*(data2[821]^data1[821])+33*(data2[820]^data1[820])+2*(data2[819]^data1[819])+2*(data2[818]^data1[818])+32*(data2[817]^data1[817])+64*(data2[816]^data1[816])+2*(data2[815]^data1[815])+2*(data2[814]^data1[814])+64*(data2[813]^data1[813])+64*(data2[812]^data1[812])+64*(data2[811]^data1[811])+64*(data2[810]^data1[810])+2*(data2[809]^data1[809])+2*(data2[808]^data1[808])+64*(data2[807]^data1[807])+2*(data2[806]^data1[806])+2*(data2[805]^data1[805])+2*(data2[804]^data1[804])+2*(data2[803]^data1[803])+33*(data2[802]^data1[802])+32*(data2[801]^data1[801])+2*(data2[800]^data1[800])+2*(data2[799]^data1[799])+2*(data2[798]^data1[798])+2*(data2[797]^data1[797])+16*(data2[796]^data1[796])+64*(data2[795]^data1[795])+2*(data2[794]^data1[794])+2*(data2[793]^data1[793])+64*(data2[792]^data1[792])+32*(data2[791]^data1[791])+2*(data2[790]^data1[790])+32*(data2[789]^data1[789])+2*(data2[788]^data1[788])+64*(data2[787]^data1[787])+64*(data2[786]^data1[786])+2*(data2[785]^data1[785])+2*(data2[784]^data1[784])+64*(data2[783]^data1[783])+64*(data2[782]^data1[782])+64*(data2[781]^data1[781])+64*(data2[780]^data1[780])+2*(data2[779]^data1[779])+2*(data2[778]^data1[778])+2*(data2[777]^data1[777])+32*(data2[776]^data1[776])+32*(data2[775]^data1[775])+64*(data2[774]^data1[774])+2*(data2[773]^data1[773])+2*(data2[772]^data1[772])+32*(data2[771]^data1[771])+32*(data2[770]^data1[770])+64*(data2[769]^data1[769])+64*(data2[768]^data1[768])+64*(data2[767]^data1[767])+2*(data2[766]^data1[766])+64*(data2[765]^data1[765])+64*(data2[764]^data1[764])+33*(data2[763]^data1[763])+64*(data2[762]^data1[762])+33*(data2[761]^data1[761])+64*(data2[760]^data1[760])+2*(data2[759]^data1[759])+32*(data2[758]^data1[758])+64*(data2[757]^data1[757])+32*(data2[756]^data1[756])+2*(data2[755]^data1[755])+64*(data2[754]^data1[754])+2*(data2[753]^data1[753])+64*(data2[752]^data1[752])+32*(data2[751]^data1[751])+2*(data2[750]^data1[750])+16*(data2[749]^data1[749])+2*(data2[748]^data1[748])+2*(data2[747]^data1[747])+16*(data2[746]^data1[746])+32*(data2[745]^data1[745])+64*(data2[744]^data1[744])+2*(data2[743]^data1[743])+32*(data2[742]^data1[742])+2*(data2[741]^data1[741])+64*(data2[740]^data1[740])+33*(data2[739]^data1[739])+2*(data2[738]^data1[738])+2*(data2[737]^data1[737])+64*(data2[736]^data1[736])+64*(data2[735]^data1[735])+33*(data2[734]^data1[734])+2*(data2[733]^data1[733])+2*(data2[732]^data1[732])+2*(data2[731]^data1[731])+64*(data2[730]^data1[730])+2*(data2[729]^data1[729])+2*(data2[728]^data1[728])+64*(data2[727]^data1[727])+64*(data2[726]^data1[726])+16*(data2[725]^data1[725])+2*(data2[724]^data1[724])+32*(data2[723]^data1[723])+32*(data2[722]^data1[722])+64*(data2[721]^data1[721])+64*(data2[720]^data1[720])+64*(data2[719]^data1[719])+2*(data2[718]^data1[718])+2*(data2[717]^data1[717])+2*(data2[716]^data1[716])+2*(data2[715]^data1[715])+2*(data2[714]^data1[714])+64*(data2[713]^data1[713])+2*(data2[712]^data1[712])+2*(data2[711]^data1[711])+64*(data2[710]^data1[710])+2*(data2[709]^data1[709])+2*(data2[708]^data1[708])+2*(data2[707]^data1[707])+64*(data2[706]^data1[706])+2*(data2[705]^data1[705])+32*(data2[704]^data1[704])+2*(data2[703]^data1[703])+64*(data2[702]^data1[702])+33*(data2[701]^data1[701])+2*(data2[700]^data1[700])+2*(data2[699]^data1[699])+64*(data2[698]^data1[698])+17*(data2[697]^data1[697])+2*(data2[696]^data1[696])+32*(data2[695]^data1[695])+32*(data2[694]^data1[694])+16*(data2[693]^data1[693])+64*(data2[692]^data1[692])+32*(data2[691]^data1[691])+64*(data2[690]^data1[690])+2*(data2[689]^data1[689])+2*(data2[688]^data1[688])+33*(data2[687]^data1[687])+2*(data2[686]^data1[686])+64*(data2[685]^data1[685])+64*(data2[684]^data1[684])+2*(data2[683]^data1[683])+64*(data2[682]^data1[682])+64*(data2[681]^data1[681])+2*(data2[680]^data1[680])+2*(data2[679]^data1[679])+2*(data2[678]^data1[678])+33*(data2[677]^data1[677])+16*(data2[676]^data1[676])+2*(data2[675]^data1[675])+64*(data2[674]^data1[674])+2*(data2[673]^data1[673])+2*(data2[672]^data1[672])+64*(data2[671]^data1[671])+2*(data2[670]^data1[670])+2*(data2[669]^data1[669])+2*(data2[668]^data1[668])+2*(data2[667]^data1[667])+2*(data2[666]^data1[666])+64*(data2[665]^data1[665])+64*(data2[664]^data1[664])+64*(data2[663]^data1[663])+64*(data2[662]^data1[662])+33*(data2[661]^data1[661])+64*(data2[660]^data1[660])+32*(data2[659]^data1[659])+64*(data2[658]^data1[658])+8*(data2[657]^data1[657])+64*(data2[656]^data1[656])+64*(data2[655]^data1[655])+2*(data2[654]^data1[654])+2*(data2[653]^data1[653])+2*(data2[652]^data1[652])+2*(data2[651]^data1[651])+2*(data2[650]^data1[650])+33*(data2[649]^data1[649])+2*(data2[648]^data1[648])+2*(data2[647]^data1[647])+64*(data2[646]^data1[646])+2*(data2[645]^data1[645])+2*(data2[644]^data1[644])+32*(data2[643]^data1[643])+2*(data2[642]^data1[642])+32*(data2[641]^data1[641])+2*(data2[640]^data1[640])+2*(data2[639]^data1[639])+2*(data2[638]^data1[638])+2*(data2[637]^data1[637])+64*(data2[636]^data1[636])+64*(data2[635]^data1[635])+64*(data2[634]^data1[634])+2*(data2[633]^data1[633])+64*(data2[632]^data1[632])+2*(data2[631]^data1[631])+2*(data2[630]^data1[630])+2*(data2[629]^data1[629])+2*(data2[628]^data1[628])+2*(data2[627]^data1[627])+33*(data2[626]^data1[626])+64*(data2[625]^data1[625])+64*(data2[624]^data1[624])+8*(data2[623]^data1[623])+64*(data2[622]^data1[622])+64*(data2[621]^data1[621])+2*(data2[620]^data1[620])+2*(data2[619]^data1[619])+33*(data2[618]^data1[618])+2*(data2[617]^data1[617])+2*(data2[616]^data1[616])+64*(data2[615]^data1[615])+32*(data2[614]^data1[614])+2*(data2[613]^data1[613])+2*(data2[612]^data1[612])+2*(data2[611]^data1[611])+2*(data2[610]^data1[610])+16*(data2[609]^data1[609])+2*(data2[608]^data1[608])+2*(data2[607]^data1[607])+64*(data2[606]^data1[606])+2*(data2[605]^data1[605])+64*(data2[604]^data1[604])+33*(data2[603]^data1[603])+2*(data2[602]^data1[602])+17*(data2[601]^data1[601])+2*(data2[600]^data1[600])+32*(data2[599]^data1[599])+32*(data2[598]^data1[598])+64*(data2[597]^data1[597])+64*(data2[596]^data1[596])+64*(data2[595]^data1[595])+64*(data2[594]^data1[594])+64*(data2[593]^data1[593])+32*(data2[592]^data1[592])+64*(data2[591]^data1[591])+2*(data2[590]^data1[590])+64*(data2[589]^data1[589])+16*(data2[588]^data1[588])+64*(data2[587]^data1[587])+9*(data2[586]^data1[586])+64*(data2[585]^data1[585])+64*(data2[584]^data1[584])+9*(data2[583]^data1[583])+2*(data2[582]^data1[582])+64*(data2[581]^data1[581])+2*(data2[580]^data1[580])+2*(data2[579]^data1[579])+64*(data2[578]^data1[578])+16*(data2[577]^data1[577])+2*(data2[576]^data1[576])+2*(data2[575]^data1[575])+2*(data2[574]^data1[574])+32*(data2[573]^data1[573])+64*(data2[572]^data1[572])+64*(data2[571]^data1[571])+32*(data2[570]^data1[570])+2*(data2[569]^data1[569])+2*(data2[568]^data1[568])+32*(data2[567]^data1[567])+33*(data2[566]^data1[566])+33*(data2[565]^data1[565])+64*(data2[564]^data1[564])+8*(data2[563]^data1[563])+64*(data2[562]^data1[562])+16*(data2[561]^data1[561])+2*(data2[560]^data1[560])+64*(data2[559]^data1[559])+2*(data2[558]^data1[558])+32*(data2[557]^data1[557])+64*(data2[556]^data1[556])+2*(data2[555]^data1[555])+2*(data2[554]^data1[554])+64*(data2[553]^data1[553])+2*(data2[552]^data1[552])+32*(data2[551]^data1[551])+64*(data2[550]^data1[550])+17*(data2[549]^data1[549])+2*(data2[548]^data1[548])+32*(data2[547]^data1[547])+64*(data2[546]^data1[546])+2*(data2[545]^data1[545])+2*(data2[544]^data1[544])+32*(data2[543]^data1[543])+64*(data2[542]^data1[542])+2*(data2[541]^data1[541])+2*(data2[540]^data1[540])+33*(data2[539]^data1[539])+2*(data2[538]^data1[538])+2*(data2[537]^data1[537])+2*(data2[536]^data1[536])+64*(data2[535]^data1[535])+33*(data2[534]^data1[534])+64*(data2[533]^data1[533])+64*(data2[532]^data1[532])+32*(data2[531]^data1[531])+32*(data2[530]^data1[530])+64*(data2[529]^data1[529])+2*(data2[528]^data1[528])+2*(data2[527]^data1[527])+2*(data2[526]^data1[526])+2*(data2[525]^data1[525])+16*(data2[524]^data1[524])+64*(data2[523]^data1[523])+2*(data2[522]^data1[522])+2*(data2[521]^data1[521])+32*(data2[520]^data1[520])+2*(data2[519]^data1[519])+32*(data2[518]^data1[518])+33*(data2[517]^data1[517])+64*(data2[516]^data1[516])+33*(data2[515]^data1[515])+16*(data2[514]^data1[514])+2*(data2[513]^data1[513])+2*(data2[512]^data1[512])+2*(data2[511]^data1[511])+2*(data2[510]^data1[510])+64*(data2[509]^data1[509])+2*(data2[508]^data1[508])+2*(data2[507]^data1[507])+2*(data2[506]^data1[506])+2*(data2[505]^data1[505])+2*(data2[504]^data1[504])+64*(data2[503]^data1[503])+64*(data2[502]^data1[502])+2*(data2[501]^data1[501])+2*(data2[500]^data1[500])+9*(data2[499]^data1[499])+2*(data2[498]^data1[498])+2*(data2[497]^data1[497])+32*(data2[496]^data1[496])+64*(data2[495]^data1[495])+64*(data2[494]^data1[494])+64*(data2[493]^data1[493])+2*(data2[492]^data1[492])+64*(data2[491]^data1[491])+2*(data2[490]^data1[490])+2*(data2[489]^data1[489])+2*(data2[488]^data1[488])+2*(data2[487]^data1[487])+16*(data2[486]^data1[486])+64*(data2[485]^data1[485])+16*(data2[484]^data1[484])+32*(data2[483]^data1[483])+2*(data2[482]^data1[482])+2*(data2[481]^data1[481])+2*(data2[480]^data1[480])+64*(data2[479]^data1[479])+2*(data2[478]^data1[478])+64*(data2[477]^data1[477])+64*(data2[476]^data1[476])+2*(data2[475]^data1[475])+33*(data2[474]^data1[474])+32*(data2[473]^data1[473])+32*(data2[472]^data1[472])+64*(data2[471]^data1[471])+64*(data2[470]^data1[470])+2*(data2[469]^data1[469])+32*(data2[468]^data1[468])+64*(data2[467]^data1[467])+64*(data2[466]^data1[466])+2*(data2[465]^data1[465])+2*(data2[464]^data1[464])+33*(data2[463]^data1[463])+2*(data2[462]^data1[462])+2*(data2[461]^data1[461])+2*(data2[460]^data1[460])+2*(data2[459]^data1[459])+64*(data2[458]^data1[458])+64*(data2[457]^data1[457])+2*(data2[456]^data1[456])+64*(data2[455]^data1[455])+2*(data2[454]^data1[454])+64*(data2[453]^data1[453])+64*(data2[452]^data1[452])+33*(data2[451]^data1[451])+2*(data2[450]^data1[450])+64*(data2[449]^data1[449])+2*(data2[448]^data1[448])+2*(data2[447]^data1[447])+64*(data2[446]^data1[446])+32*(data2[445]^data1[445])+64*(data2[444]^data1[444])+2*(data2[443]^data1[443])+2*(data2[442]^data1[442])+2*(data2[441]^data1[441])+2*(data2[440]^data1[440])+2*(data2[439]^data1[439])+64*(data2[438]^data1[438])+2*(data2[437]^data1[437])+2*(data2[436]^data1[436])+32*(data2[435]^data1[435])+64*(data2[434]^data1[434])+2*(data2[433]^data1[433])+64*(data2[432]^data1[432])+33*(data2[431]^data1[431])+64*(data2[430]^data1[430])+2*(data2[429]^data1[429])+32*(data2[428]^data1[428])+32*(data2[427]^data1[427])+64*(data2[426]^data1[426])+2*(data2[425]^data1[425])+33*(data2[424]^data1[424])+64*(data2[423]^data1[423])+64*(data2[422]^data1[422])+2*(data2[421]^data1[421])+2*(data2[420]^data1[420])+2*(data2[419]^data1[419])+2*(data2[418]^data1[418])+64*(data2[417]^data1[417])+33*(data2[416]^data1[416])+2*(data2[415]^data1[415])+64*(data2[414]^data1[414])+2*(data2[413]^data1[413])+32*(data2[412]^data1[412])+32*(data2[411]^data1[411])+32*(data2[410]^data1[410])+64*(data2[409]^data1[409])+2*(data2[408]^data1[408])+64*(data2[407]^data1[407])+2*(data2[406]^data1[406])+64*(data2[405]^data1[405])+64*(data2[404]^data1[404])+2*(data2[403]^data1[403])+2*(data2[402]^data1[402])+33*(data2[401]^data1[401])+2*(data2[400]^data1[400])+8*(data2[399]^data1[399])+64*(data2[398]^data1[398])+2*(data2[397]^data1[397])+64*(data2[396]^data1[396])+64*(data2[395]^data1[395])+2*(data2[394]^data1[394])+8*(data2[393]^data1[393])+33*(data2[392]^data1[392])+32*(data2[391]^data1[391])+2*(data2[390]^data1[390])+32*(data2[389]^data1[389])+2*(data2[388]^data1[388])+64*(data2[387]^data1[387])+64*(data2[386]^data1[386])+64*(data2[385]^data1[385])+2*(data2[384]^data1[384])+2*(data2[383]^data1[383])+64*(data2[382]^data1[382])+32*(data2[381]^data1[381])+64*(data2[380]^data1[380])+2*(data2[379]^data1[379])+64*(data2[378]^data1[378])+64*(data2[377]^data1[377])+16*(data2[376]^data1[376])+64*(data2[375]^data1[375])+2*(data2[374]^data1[374])+2*(data2[373]^data1[373])+64*(data2[372]^data1[372])+64*(data2[371]^data1[371])+64*(data2[370]^data1[370])+2*(data2[369]^data1[369])+2*(data2[368]^data1[368])+2*(data2[367]^data1[367])+2*(data2[366]^data1[366])+2*(data2[365]^data1[365])+2*(data2[364]^data1[364])+33*(data2[363]^data1[363])+16*(data2[362]^data1[362])+64*(data2[361]^data1[361])+2*(data2[360]^data1[360])+2*(data2[359]^data1[359])+2*(data2[358]^data1[358])+2*(data2[357]^data1[357])+64*(data2[356]^data1[356])+64*(data2[355]^data1[355])+64*(data2[354]^data1[354])+2*(data2[353]^data1[353])+2*(data2[352]^data1[352])+32*(data2[351]^data1[351])+16*(data2[350]^data1[350])+2*(data2[349]^data1[349])+32*(data2[348]^data1[348])+2*(data2[347]^data1[347])+2*(data2[346]^data1[346])+8*(data2[345]^data1[345])+16*(data2[344]^data1[344])+33*(data2[343]^data1[343])+16*(data2[342]^data1[342])+2*(data2[341]^data1[341])+64*(data2[340]^data1[340])+16*(data2[339]^data1[339])+2*(data2[338]^data1[338])+8*(data2[337]^data1[337])+64*(data2[336]^data1[336])+64*(data2[335]^data1[335])+2*(data2[334]^data1[334])+2*(data2[333]^data1[333])+2*(data2[332]^data1[332])+32*(data2[331]^data1[331])+2*(data2[330]^data1[330])+2*(data2[329]^data1[329])+64*(data2[328]^data1[328])+16*(data2[327]^data1[327])+2*(data2[326]^data1[326])+2*(data2[325]^data1[325])+2*(data2[324]^data1[324])+2*(data2[323]^data1[323])+16*(data2[322]^data1[322])+2*(data2[321]^data1[321])+32*(data2[320]^data1[320])+64*(data2[319]^data1[319])+16*(data2[318]^data1[318])+2*(data2[317]^data1[317])+32*(data2[316]^data1[316])+2*(data2[315]^data1[315])+64*(data2[314]^data1[314])+16*(data2[313]^data1[313])+2*(data2[312]^data1[312])+32*(data2[311]^data1[311])+32*(data2[310]^data1[310])+64*(data2[309]^data1[309])+64*(data2[308]^data1[308])+2*(data2[307]^data1[307])+2*(data2[306]^data1[306])+32*(data2[305]^data1[305])+33*(data2[304]^data1[304])+2*(data2[303]^data1[303])+32*(data2[302]^data1[302])+2*(data2[301]^data1[301])+17*(data2[300]^data1[300])+64*(data2[299]^data1[299])+2*(data2[298]^data1[298])+64*(data2[297]^data1[297])+2*(data2[296]^data1[296])+2*(data2[295]^data1[295])+64*(data2[294]^data1[294])+64*(data2[293]^data1[293])+32*(data2[292]^data1[292])+32*(data2[291]^data1[291])+2*(data2[290]^data1[290])+64*(data2[289]^data1[289])+64*(data2[288]^data1[288])+2*(data2[287]^data1[287])+2*(data2[286]^data1[286])+64*(data2[285]^data1[285])+64*(data2[284]^data1[284])+2*(data2[283]^data1[283])+32*(data2[282]^data1[282])+32*(data2[281]^data1[281])+2*(data2[280]^data1[280])+2*(data2[279]^data1[279])+2*(data2[278]^data1[278])+2*(data2[277]^data1[277])+16*(data2[276]^data1[276])+32*(data2[275]^data1[275])+9*(data2[274]^data1[274])+9*(data2[273]^data1[273])+64*(data2[272]^data1[272])+32*(data2[271]^data1[271])+2*(data2[270]^data1[270])+2*(data2[269]^data1[269])+2*(data2[268]^data1[268])+64*(data2[267]^data1[267])+33*(data2[266]^data1[266])+2*(data2[265]^data1[265])+2*(data2[264]^data1[264])+2*(data2[263]^data1[263])+64*(data2[262]^data1[262])+64*(data2[261]^data1[261])+2*(data2[260]^data1[260])+16*(data2[259]^data1[259])+32*(data2[258]^data1[258])+32*(data2[257]^data1[257])+32*(data2[256]^data1[256])+16*(data2[255]^data1[255])+2*(data2[254]^data1[254])+64*(data2[253]^data1[253])+32*(data2[252]^data1[252])+64*(data2[251]^data1[251])+2*(data2[250]^data1[250])+2*(data2[249]^data1[249])+2*(data2[248]^data1[248])+2*(data2[247]^data1[247])+32*(data2[246]^data1[246])+64*(data2[245]^data1[245])+64*(data2[244]^data1[244])+2*(data2[243]^data1[243])+2*(data2[242]^data1[242])+2*(data2[241]^data1[241])+2*(data2[240]^data1[240])+64*(data2[239]^data1[239])+2*(data2[238]^data1[238])+2*(data2[237]^data1[237])+2*(data2[236]^data1[236])+32*(data2[235]^data1[235])+2*(data2[234]^data1[234])+64*(data2[233]^data1[233])+8*(data2[232]^data1[232])+2*(data2[231]^data1[231])+2*(data2[230]^data1[230])+2*(data2[229]^data1[229])+64*(data2[228]^data1[228])+64*(data2[227]^data1[227])+64*(data2[226]^data1[226])+33*(data2[225]^data1[225])+2*(data2[224]^data1[224])+16*(data2[223]^data1[223])+2*(data2[222]^data1[222])+2*(data2[221]^data1[221])+16*(data2[220]^data1[220])+2*(data2[219]^data1[219])+2*(data2[218]^data1[218])+64*(data2[217]^data1[217])+2*(data2[216]^data1[216])+33*(data2[215]^data1[215])+64*(data2[214]^data1[214])+2*(data2[213]^data1[213])+64*(data2[212]^data1[212])+2*(data2[211]^data1[211])+2*(data2[210]^data1[210])+8*(data2[209]^data1[209])+64*(data2[208]^data1[208])+64*(data2[207]^data1[207])+2*(data2[206]^data1[206])+2*(data2[205]^data1[205])+2*(data2[204]^data1[204])+64*(data2[203]^data1[203])+64*(data2[202]^data1[202])+2*(data2[201]^data1[201])+2*(data2[200]^data1[200])+2*(data2[199]^data1[199])+32*(data2[198]^data1[198])+2*(data2[197]^data1[197])+16*(data2[196]^data1[196])+2*(data2[195]^data1[195])+2*(data2[194]^data1[194])+64*(data2[193]^data1[193])+2*(data2[192]^data1[192])+64*(data2[191]^data1[191])+64*(data2[190]^data1[190])+16*(data2[189]^data1[189])+64*(data2[188]^data1[188])+2*(data2[187]^data1[187])+64*(data2[186]^data1[186])+64*(data2[185]^data1[185])+64*(data2[184]^data1[184])+64*(data2[183]^data1[183])+2*(data2[182]^data1[182])+33*(data2[181]^data1[181])+2*(data2[180]^data1[180])+2*(data2[179]^data1[179])+32*(data2[178]^data1[178])+2*(data2[177]^data1[177])+32*(data2[176]^data1[176])+2*(data2[175]^data1[175])+64*(data2[174]^data1[174])+64*(data2[173]^data1[173])+2*(data2[172]^data1[172])+2*(data2[171]^data1[171])+33*(data2[170]^data1[170])+2*(data2[169]^data1[169])+16*(data2[168]^data1[168])+64*(data2[167]^data1[167])+2*(data2[166]^data1[166])+2*(data2[165]^data1[165])+2*(data2[164]^data1[164])+64*(data2[163]^data1[163])+2*(data2[162]^data1[162])+2*(data2[161]^data1[161])+2*(data2[160]^data1[160])+2*(data2[159]^data1[159])+64*(data2[158]^data1[158])+64*(data2[157]^data1[157])+64*(data2[156]^data1[156])+2*(data2[155]^data1[155])+2*(data2[154]^data1[154])+2*(data2[153]^data1[153])+2*(data2[152]^data1[152])+2*(data2[151]^data1[151])+2*(data2[150]^data1[150])+64*(data2[149]^data1[149])+2*(data2[148]^data1[148])+64*(data2[147]^data1[147])+32*(data2[146]^data1[146])+8*(data2[145]^data1[145])+16*(data2[144]^data1[144])+33*(data2[143]^data1[143])+32*(data2[142]^data1[142])+32*(data2[141]^data1[141])+2*(data2[140]^data1[140])+2*(data2[139]^data1[139])+32*(data2[138]^data1[138])+32*(data2[137]^data1[137])+2*(data2[136]^data1[136])+64*(data2[135]^data1[135])+9*(data2[134]^data1[134])+2*(data2[133]^data1[133])+2*(data2[132]^data1[132])+32*(data2[131]^data1[131])+16*(data2[130]^data1[130])+2*(data2[129]^data1[129])+2*(data2[128]^data1[128])+32*(data2[127]^data1[127])+32*(data2[126]^data1[126])+2*(data2[125]^data1[125])+64*(data2[124]^data1[124])+32*(data2[123]^data1[123])+2*(data2[122]^data1[122])+16*(data2[121]^data1[121])+64*(data2[120]^data1[120])+2*(data2[119]^data1[119])+2*(data2[118]^data1[118])+2*(data2[117]^data1[117])+16*(data2[116]^data1[116])+2*(data2[115]^data1[115])+2*(data2[114]^data1[114])+16*(data2[113]^data1[113])+64*(data2[112]^data1[112])+32*(data2[111]^data1[111])+2*(data2[110]^data1[110])+64*(data2[109]^data1[109])+33*(data2[108]^data1[108])+2*(data2[107]^data1[107])+2*(data2[106]^data1[106])+64*(data2[105]^data1[105])+2*(data2[104]^data1[104])+64*(data2[103]^data1[103])+32*(data2[102]^data1[102])+32*(data2[101]^data1[101])+64*(data2[100]^data1[100])+33*(data2[99]^data1[99])+2*(data2[98]^data1[98])+2*(data2[97]^data1[97])+64*(data2[96]^data1[96])+64*(data2[95]^data1[95])+64*(data2[94]^data1[94])+2*(data2[93]^data1[93])+32*(data2[92]^data1[92])+9*(data2[91]^data1[91])+32*(data2[90]^data1[90])+2*(data2[89]^data1[89])+64*(data2[88]^data1[88])+64*(data2[87]^data1[87])+2*(data2[86]^data1[86])+64*(data2[85]^data1[85])+64*(data2[84]^data1[84])+2*(data2[83]^data1[83])+2*(data2[82]^data1[82])+2*(data2[81]^data1[81])+2*(data2[80]^data1[80])+2*(data2[79]^data1[79])+16*(data2[78]^data1[78])+2*(data2[77]^data1[77])+64*(data2[76]^data1[76])+2*(data2[75]^data1[75])+64*(data2[74]^data1[74])+2*(data2[73]^data1[73])+2*(data2[72]^data1[72])+32*(data2[71]^data1[71])+64*(data2[70]^data1[70])+64*(data2[69]^data1[69])+64*(data2[68]^data1[68])+2*(data2[67]^data1[67])+2*(data2[66]^data1[66])+2*(data2[65]^data1[65])+32*(data2[64]^data1[64])+2*(data2[63]^data1[63])+2*(data2[62]^data1[62])+64*(data2[61]^data1[61])+64*(data2[60]^data1[60])+64*(data2[59]^data1[59])+2*(data2[58]^data1[58])+64*(data2[57]^data1[57])+16*(data2[56]^data1[56])+2*(data2[55]^data1[55])+2*(data2[54]^data1[54])+16*(data2[53]^data1[53])+64*(data2[52]^data1[52])+64*(data2[51]^data1[51])+2*(data2[50]^data1[50])+16*(data2[49]^data1[49])+64*(data2[48]^data1[48])+17*(data2[47]^data1[47])+2*(data2[46]^data1[46])+2*(data2[45]^data1[45])+2*(data2[44]^data1[44])+32*(data2[43]^data1[43])+16*(data2[42]^data1[42])+32*(data2[41]^data1[41])+64*(data2[40]^data1[40])+2*(data2[39]^data1[39])+2*(data2[38]^data1[38])+64*(data2[37]^data1[37])+64*(data2[36]^data1[36])+64*(data2[35]^data1[35])+32*(data2[34]^data1[34])+2*(data2[33]^data1[33])+33*(data2[32]^data1[32])+2*(data2[31]^data1[31])+2*(data2[30]^data1[30])+2*(data2[29]^data1[29])+64*(data2[28]^data1[28])+64*(data2[27]^data1[27])+2*(data2[26]^data1[26])+2*(data2[25]^data1[25])+2*(data2[24]^data1[24])+2*(data2[23]^data1[23])+2*(data2[22]^data1[22])+64*(data2[21]^data1[21])+32*(data2[20]^data1[20])+32*(data2[19]^data1[19])+16*(data2[18]^data1[18])+64*(data2[17]^data1[17])+2*(data2[16]^data1[16])+2*(data2[15]^data1[15])+64*(data2[14]^data1[14])+16*(data2[13]^data1[13])+17*(data2[12]^data1[12])+64*(data2[11]^data1[11])+2*(data2[10]^data1[10])+32*(data2[9]^data1[9])+64*(data2[8]^data1[8])+2*(data2[7]^data1[7])+16*(data2[6]^data1[6])+2*(data2[5]^data1[5])+64*(data2[4]^data1[4])+2*(data2[3]^data1[3])+33*(data2[2]^data1[2])+64*(data2[1]^data1[1])+64*(data2[0]^data1[0]));
		end
		integer w_file;
		initial w_file = $fopen("semifixed_L_trace.txt", "w");
always @(posedge clk)
    begin
        //$fdisplay(w_file,"%d",trig);
        $fwrite(w_file,"%d\n",$signed(plot));
    end	 


      
endmodule

